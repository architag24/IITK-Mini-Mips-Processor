module instruction_mem (
    input [31:0] addr,
    output [31:0] instruction
);
    reg [31:0] memory [0:255]; // 1 KB instr mem
//    memory[31] =

    initial begin

        //insertion sort

         memory[0] = 32'b00100000000111110000000000000111;  //storing number of values=7 for insertion sort in $31
         memory[1] = 32'b00100000000000010000000000000000; // addi $1, $0, 0
         memory[2] = 32'b00100000001000010000000000000001; // addi $1, $1, 1
         memory[3] = 32'b00010000001111110000000001100100; // beq  $1, $31, 100
         memory[4] = 32'b00100000001000101111111111111111; // addi $2, $1, -1
         memory[5] = 32'b00100000010001010000000000000001; // add  $5, $2, 1
         memory[6] = 32'b10001100010001110000000000000000; // lw   $7, 0($2)
         memory[7] = 32'b10001100101010000000000000000000; // lw   $8, 0($5)
         memory[8] = 32'b00010100111010001111111111111001; // bleq $7, $8, -7
         memory[9] = 32'b10101100101001110000000000000000; // sw   $7, 0($5)
         memory[10] = 32'b10101100010010000000000000000000; // sw   $8, 0($2)
         memory[11] = 32'b00010000010000001111111111110110; // beq  $2, $0, -10
         memory[12] = 32'b00100000010000101111111111111111; // addi $2, $2, -1
         memory[13] = 32'b00010000000000001111111111110111; // beq  $0, $0, -9
//         memory[0] = 32'b00100000000010000000000000001010; // addi $8, $0, 10
//         memory[1] = 32'b00100000000010010000000000000110; // addi $9, $0, 6
//         memory[2] = 32'b00010101000010010000000000000010; // bleq  $8, $9, label (offset = 2)
//         memory[3] = 32'b00100000000010100000000011111111; // addi $10, $0, 255 (skipped if branch taken)
//         memory[4] = 32'b00100000000010110000000000001010; // addi $11, $0, 10
//         memory[5] = 32'b00000001000010010110000000011000; // mul-low $12, $8, $9
         //memory[6] = 32'b00000001000010            // mul-high $13 ,$8,$9

//         memory[0] = 32'b00100000000010000000000000000101; // addi $8, $0, 5
//         memory[1] = 32'b00100000000010010000000000001010; // addi $9, $0, 10
//         memory[2] = 32'b00000001000010010101000000100000; // add  $10,$8,$9
//         memory[3] = 32'b10101101000010100000000000000000; // sw   $10, 0($8)
//         memory[4] = 32'b10001101000010110000000000000000; // lw   $11, 0($8)

    end

    assign instruction = memory[addr[31:2]]; // word-aligned
endmodule

